
`timescale 1 ns / 1 ps

module axis_master_data_gen_mem#
(
    parameter integer C_M_AXIS_TDATA_WIDTH	= 32,
    parameter integer C_M_START_COUNT	= 32
)
(
    m00_axis_aclk,
    m00_axis_aresetn,
    m00_axis_tvalid,
    m00_axis_tdata,
    m00_axis_tstrb,
    m00_axis_tlast,
    m00_axis_tready
);
    input                                              m00_axis_aclk;
    input                                              m00_axis_aresetn;
    output                                             m00_axis_tvalid;
    output   [C_M_AXIS_TDATA_WIDTH-1 : 0]              m00_axis_tdata;
    output   [(C_M_AXIS_TDATA_WIDTH/8)-1 : 0]          m00_axis_tstrb;
    output                                             m00_axis_tlast;
    input                                              m00_axis_tready;

    /*
        User controlled parameters
    */
    // localparam NUMBER_OF_OUTPUT_WORDS = 100;//261;
    localparam NUMBER_OF_OUTPUT_WORDS = 20;//261;
    localparam OUTPUT_WORD_ID_STALL_FOR_50_CYCLE = NUMBER_OF_OUTPUT_WORDS-4;//261;

    function integer clogb2 (input integer bit_depth);
        begin
            for(clogb2=0; bit_depth>0; clogb2=clogb2+1)
                bit_depth = bit_depth >> 1;
        end
    endfunction

    reg [$clog2(NUMBER_OF_OUTPUT_WORDS)-1:0]           read_pointer;
    reg [C_M_AXIS_TDATA_WIDTH-1:0]                     m00_axis_tdata_inner;
    reg                                                m00_axis_tvalid_inner;
    wire                                               send_tx;
    assign    send_tx = m00_axis_tvalid_inner & m00_axis_tready;
    reg                                                tx_done;
    reg                                                no_send;
    reg      [$clog2(NUMBER_OF_OUTPUT_WORDS)-1:0]      stall_cnt;

    reg      [C_M_AXIS_TDATA_WIDTH-1:0]                mem[0:NUMBER_OF_OUTPUT_WORDS-1];
    initial
    begin
        stall_cnt <= 0;
        mem[0] = 128'b00000000000000000000000000000000000000000000000000000000111010001111100010111010111111001001111101110111110000111110110000100001;
        mem[1] = 128'b00000000000000000000000000000000000000000000000000000000111100110001011001111000010111110010001001110111110010111111101000001110;
        mem[2] = 128'b00000000000000000000000000000000000000000000000000000000000011101000001001000101011000100100000000100000000110000001011111110010;
        mem[3] = 128'b00000000000000000000000000000000000000000000000000000000001001100111101000111100011000101001111110100000000101111111101111111101;
        mem[4] = 128'b00000000000000000000000000000000000000000000000000000000001111001001111010111110000001111111000101110111001110001100000000101001;
        mem[5] = 128'b00000000000000000000000000000000000000000000000000000000000111011111100111000101001000101001000000100000010010000100111111101100;
        mem[6] = 128'b00000000000000000000000000000000000000000000000000000000110110110000010101000011001111011110000001010111111011000000111111111111;
        mem[7] = 128'b00000000000000000000000000000000000000000000000000000000111001111111111100111101010111101110111111011001010100001000011000001001;
        mem[8] = 128'b00000000000000000000000000000000000000000000000000000000111101010111100101111101111111101011111101010111101101111101011111101101;
        mem[9] = 128'b00000000000000000000000000000000000000000000000000000000111110101111101111111110110111110010111101111111110100111110000111101101;
        mem[10] = 128'b00000000000000000000000000000000000000000000000000000000111111000111110110111110011111111000111110110111110100111110111111110100;
        mem[11] = 128'b00000000000000000000000000000000000000000000000000000000111101111111110100111101011111101111111110011111101011111101111111110100;
        mem[12] = 128'b00000000000000000000000000000000000000000000000000000000111101111111101101111110001111101101111101011111110010111101110111101011;
        mem[13] = 128'b00000000000000000000000000000000000000000000000000000000111110110111110011111110111111110101111110001111110111111110100111110010;
        mem[14] = 128'b00000000000000000000000000000000000000000000000000000000111110100111111000111101111111110010111110111111101110111110010111110111;
        mem[15] = 128'b00000000000000000000000000000000000000000000000000000000111101111111110000111110010111101110111101111111110001111101111111101110;
        // mem[0] = 128'b00000000000000000000000000000000000000000000000000000000111010001111100010111010111111001001111101110111110000111110110000100001;
        // mem[1] = 128'b00000000000000000000000000000000000000000000000000000000111100110001011001111000010111110010001001110111110010111111101000001110;
        // mem[2] = 128'b00000000000000000000000000000000000000000000000000000000000011101000001001000101011000100100000000100000000110000001011111110010;
        // mem[3] = 128'b00000000000000000000000000000000000000000000000000000000001001100111101000111100011000101001111110100000000101111111101111111101;
        // mem[4] = 128'b00000000000000000000000000000000000000000000000000000000001111001001111010111110000001111111000101110111001110001100000000101001;
        // mem[5] = 128'b00000000000000000000000000000000000000000000000000000000000111011111100111000101001000101001000000100000010010000100111111101100;
        // mem[6] = 128'b00000000000000000000000000000000000000000000000000000000110110110000010101000011001111011110000001010111111011000000111111111111;
        // mem[7] = 128'b00000000000000000000000000000000000000000000000000000000111001111111111100111101010111101110111111011001010100001000011000001001;
        // mem[8] = 128'b00000000000000000000000000000000000000000000000000000000000010000000000000000010011000010011000000000000000000000000000000000000;
        // mem[9] = 128'b00000000000000000000000000000000000000000000000000000000000001111000010000000010100000010100000010011000000000000000000000000000;
        // mem[10] = 128'b00000000000000000000000000000000000000000000000000000000000010010000010001000010101000010101000010100000000000000000000000000000;
        // mem[11] = 128'b00000000000000000000000000000000000000000000000000000000000010100000010101000010010000010100000010101000000000000000000000000000;
        // mem[12] = 128'b00000000000000000000000000000000000000000000000000000000000010110000010101000010010000010010000010010000000000000000000000000000;
        // mem[13] = 128'b00000000000000000000000000000000000000000000000000000000000011001000010111000010011000010011000010010000000000000000000000000000;
        // mem[14] = 128'b00000000000000000000000000000000000000000000000000000000000011010000011010000010110000010011000010011000000000000000000000000000;
        // mem[15] = 128'b00000000000000000000000000000000000000000000000000000000000011100000011011000011000000010111000010110000000000000000000000000000;
        // mem[16] = 128'b00000000000000000000000000000000000000000000000000000000000011100000011010000011011000011010000011000000000000000000000000000000;
        // mem[17] = 128'b00000000000000000000000000000000000000000000000000000000000011001000011010000010111000011010000011011000000000000000000000000000;
        // mem[18] = 128'b00000000000000000000000000000000000000000000000000000000000010110000011010000011001000010111000010111000000000000000000000000000;
        // mem[19] = 128'b00000000000000000000000000000000000000000000000000000000000010110000011000000010110000010111000011001000000000000000000000000000;
        // mem[20] = 128'b00000000000000000000000000000000000000000000000000000000000010110000010101000011011000011000000010110000000000000000000000000000;
        // mem[21] = 128'b00000000000000000000000000000000000000000000000000000000000011011000011001000011110000011101000011011000000000000000000000000000;
        // mem[22] = 128'b00000000000000000000000000000000000000000000000000000000000011011000011100000011011000011101000011110000000000000000000000000000;
        // mem[23] = 128'b00000000000000000000000000000000000000000000000000000000000011000000011001000011010000011100000011011000000000000000000000000000;
        // mem[24] = 128'b00000000000000000000000000000000000000000000000000000000000011001000011000000010111000011001000011010000000000000000000000000000;
        // mem[25] = 128'b00000000000000000000000000000000000000000000000000000000000010110000010111000001110000011000000010111000000000000000000000000000;
        // mem[26] = 128'b00000000000000000000000000000000000000000000000000000000000000111000010000111111101000000111000001110000000000000000000000000000;
        // mem[27] = 128'b00000000000000000000000000000000000000000000000000000000111110111111111101111110101111110111111111101000000000000000000000000000;
        // mem[28] = 128'b00000000000000000000000000000000000000000000000000000000111110001111110111111110010111110001111110101000000000000000000000000000;
        // mem[29] = 128'b00000000000000000000000000000000000000000000000000000000111110110111110010111111110111110111111110010000000000000000000000000000;
        // mem[30] = 128'b00000000000000000000000000000000000000000000000000000000111111011111111100111111001111111100111111110000000000000000000000000000;
        // mem[31] = 128'b00000000000000000000000000000000000000000000000000000000111110111111110111111111000111111000111111001000000000000000000000000000;
        // mem[32] = 128'b00000000000000000000000000000000000000000000000000000000111110111111111000111110110111110111111111000000000000000000000000000000;
        // mem[33] = 128'b00000000000000000000000000000000000000000000000000000000111111000111110101111110110111111000111110110000000000000000000000000000;
        // mem[34] = 128'b00000000000000000000000000000000000000000000000000000000111110100111110111111101101111110010111110110000000000000000000000000000;
        // mem[35] = 128'b00000000000000000000000000000000000000000000000000000000111101011111101111111101000111101001111101101000000000000000000000000000;
        // mem[36] = 128'b00000000000000000000000000000000000000000000000000000000111101001111101000111101011111101000111101000000000000000000000000000000;
        // mem[37] = 128'b00000000000000000000000000000000000000000000000000000000111101100111101011111101101111101101111101011000000000000000000000000000;
        // mem[38] = 128'b00000000000000000000000000000000000000000000000000000000111101010111101011111101010111101011111101101000000000000000000000000000;
        // mem[39] = 128'b00000000000000000000000000000000000000000000000000000000111101001111101010111100111111101010111101010000000000000000000000000000;
        // mem[40] = 128'b00000000000000000000000000000000000000000000000000000000111100011111101000111101000111100110111100111000000000000000000000000000;
        // mem[41] = 128'b00000000000000000000000000000000000000000000000000000000111101000111100111111101001111101001111101000000000000000000000000000000;
        // mem[42] = 128'b00000000000000000000000000000000000000000000000000000000111101001111101001111101000111101000111101001000000000000000000000000000;
        // mem[43] = 128'b00000000000000000000000000000000000000000000000000000000111101001111101001111101000111101000111101000000000000000000000000000000;
        // mem[44] = 128'b00000000000000000000000000000000000000000000000000000000111101000111101000111101010111101001111101000000000000000000000000000000;
        // mem[45] = 128'b00000000000000000000000000000000000000000000000000000000111100110111101010111100101111101000111101010000000000000000000000000000;
        // mem[46] = 128'b00000000000000000000000000000000000000000000000000000000111100010111100011111011110111100011111100101000000000000000000000000000;
        // mem[47] = 128'b00000000000000000000000000000000000000000000000000000000111011101111011100111011101111011110111011110000000000000000000000000000;
        // mem[48] = 128'b00000000000000000000000000000000000000000000000000000000111011110111011100111011111111011101111011101000000000000000000000000000;
        // mem[49] = 128'b00000000000000000000000000000000000000000000000000000000111100111111100010111100111111100100111011111000000000000000000000000000;
        // mem[50] = 128'b00000000000000000000000000000000000000000000000000000000111101010111101001111101000111101001111100111000000000000000000000000000;
        // mem[51] = 128'b00000000000000000000000000000000000000000000000000000000111101001111101000111101111111101011111101000000000000000000000000000000;
        // mem[52] = 128'b00000000000000000000000000000000000000000000000000000000111101100111101111111100100111101101111101111000000000000000000000000000;
        // mem[53] = 128'b00000000000000000000000000000000000000000000000000000000111011101111100101111011101111011101111100100000000000000000000000000000;
        // mem[54] = 128'b00000000000000000000000000000000000000000000000000000000111011110111011011111011111111011110111011101000000000000000000000000000;
        // mem[55] = 128'b00000000000000000000000000000000000000000000000000000000111011010111011110111010110111011010111011111000000000000000000000000000;
        // mem[56] = 128'b00000000000000000000000000000000000000000000000000000000111010101111010110111010101111010100111010110000000000000000000000000000;
        // mem[57] = 128'b00000000000000000000000000000000000000000000000000000000111010111111010110111011000111010111111010101000000000000000000000000000;
        // mem[58] = 128'b00000000000000000000000000000000000000000000000000000000111011001111010111111011101111011010111011000000000000000000000000000000;
        // mem[59] = 128'b00000000000000000000000000000000000000000000000000000000111100001111011100111100101111100011111011101000000000000000000000000000;
        // mem[60] = 128'b00000000000000000000000000000000000000000000000000000000111100101111100110111100101111100101111100101000000000000000000000000000;
        // mem[61] = 128'b00000000000000000000000000000000000000000000000000000000111100101111100101111100101111100100111100101000000000000000000000000000;
        // mem[62] = 128'b00000000000000000000000000000000000000000000000000000000111101011111100111111110001111101010111100101000000000000000000000000000;
        // mem[63] = 128'b00000000000000000000000000000000000000000000000000000000111110010111110011111101111111110000111110001000000000000000000000000000;
        // mem[64] = 128'b00000000000000000000000000000000000000000000000000000000111101100111110000111101011111101100111101111000000000000000000000000000;
        // mem[65] = 128'b00000000000000000000000000000000000000000000000000000000111101100111101010111110000111101100111101011000000000000000000000000000;
        // mem[66] = 128'b00000000000000000000000000000000000000000000000000000000111110000111110000111110010111110011111110000000000000000000000000000000;
        // mem[67] = 128'b00000000000000000000000000000000000000000000000000000000111101110111110010111101111111110000111110010000000000000000000000000000;
        // mem[68] = 128'b00000000000000000000000000000000000000000000000000000000111101111111101100111110011111110000111101111000000000000000000000000000;
        // mem[69] = 128'b00000000000000000000000000000000000000000000000000000000111110011111110010111110010111110100111110011000000000000000000000000000;
        // mem[70] = 128'b00000000000000000000000000000000000000000000000000000000111101111111110011111101101111110000111110010000000000000000000000000000;
        // mem[71] = 128'b00000000000000000000000000000000000000000000000000000000111101011111101100111101100111101100111101101000000000000000000000000000;
        // mem[72] = 128'b00000000000000000000000000000000000000000000000000000000111110001111101100111110101111110001111101100000000000000000000000000000;
        // mem[73] = 128'b00000000000000000000000000000000000000000000000000000000111111000111110101111110101111110111111110101000000000000000000000000000;
        // mem[74] = 128'b00000000000000000000000000000000000000000000000000000000111101101111110011111101010111101101111110101000000000000000000000000000;
        // mem[75] = 128'b00000000000000000000000000000000000000000000000000000000111101101111101011111110101111101101111101010000000000000000000000000000;
        // mem[76] = 128'b00000000000000000000000000000000000000000000000000000000111111000111110010111111000111111000111110101000000000000000000000000000;
        // mem[77] = 128'b00000000000000000000000000000000000000000000000000000000111110100111110111111101111111110100111111000000000000000000000000000000;
        // mem[78] = 128'b00000000000000000000000000000000000000000000000000000000111101110111110000111110011111110000111101111000000000000000000000000000;
        // mem[79] = 128'b00000000000000000000000000000000000000000000000000000000111110010111110010111101101111110011111110011000000000000000000000000000;
        // mem[80] = 128'b00000000000000000000000000000000000000000000000000000000111101111111101101111110010111101001111101101000000000000000000000000000;
        // mem[81] = 128'b00000000000000000000000000000000000000000000000000000000000001011111111110000001111000000100111110010000000000000000000000000000;
        // mem[82] = 128'b00000000000000000000000000000000000000000000000000000000000001010000001110000001001000000111000001111000000000000000000000000000;
        // mem[83] = 128'b00000000000000000000000000000000000000000000000000000000000001110000001100000001101000001110000001001000000000000000000000000000;
        // mem[84] = 128'b00000000000000000000000000000000000000000000000000000000000010010000001111000010000000001111000001101000000000000000000000000000;
        // mem[85] = 128'b00000000000000000000000000000000000000000000000000000000000010011000010011000010000000010000000010000000000000000000000000000000;
        // mem[86] = 128'b00000000000000000000000000000000000000000000000000000000000010101000010011000010100000010010000010000000000000000000000000000000;
        // mem[87] = 128'b00000000000000000000000000000000000000000000000000000000000010011000010101000010001000010100000010100000000000000000000000000000;
        // mem[88] = 128'b00000000000000000000000000000000000000000000000000000000000010001000010010000010000000001111000010001000000000000000000000000000;
        // mem[89] = 128'b00000000000000000000000000000000000000000000000000000000000001101000010001000010000000010000000010000000000000000000000000000000;
        // mem[90] = 128'b00000000000000000000000000000000000000000000000000000000000010000000001011000001111000001100000010000000000000000000000000000000;
        // mem[91] = 128'b00000000000000000000000000000000000000000000000000000000000010110000010011000010100000010010000001111000000000000000000000000000;
        // mem[92] = 128'b00000000000000000000000000000000000000000000000000000000000011100000011011000010110000010011000010100000000000000000000000000000;
        // mem[93] = 128'b00000000000000000000000000000000000000000000000000000000000101111000100010000111000000100111000010110000000000000000000000000000;
        // mem[94] = 128'b00000000000000000000000000000000000000000000000000000000000111001000111010000111011000111011000111000000000000000000000000000000;
        // mem[95] = 128'b00000000000000000000000000000000000000000000000000000000000100111000110001000110101000111001000111011000000000000000000000000000;
        // mem[96] = 128'b00000000000000000000000000000000000000000000000000000000000011010000011111000100010000101011000110101000000000000000000000000000;
        // mem[97] = 128'b00000000000000000000000000000000000000000000000000000000000010011000010101000010101000011010000100010000000000000000000000000000;
        // mem[98] = 128'b00000000000000000000000000000000000000000000000000000000000010001000010001000010010000010110000010101000000000000000000000000000;
        // mem[99] = 128'b00000000000000000000000000000000000000000000000000000000000010001000010001000001110000001101000010010000000000000000000000000000;
        // mem[100] = 128'b00000000000000000000000000000000000000000000000000000000000001101000001110000001100000001101000001110000000000000000000000000000;
        // mem[101] = 128'b00000000000000000000000000000000000000000000000000000000000001100000001101000001010000001010000001100000000000000000000000000000;
        // mem[102] = 128'b00000000000000000000000000000000000000000000000000000000000010011000001111000010001000001101000001010000000000000000000000000000;
        // mem[103] = 128'b00000000000000000000000000000000000000000000000000000000000010000000010100000000111000010001000010001000000000000000000000000000;
        // mem[104] = 128'b00000000000000000000000000000000000000000000000000000000111111101000000101111111110000000001000000111000000000000000000000000000;
        // mem[105] = 128'b00000000000000000000000000000000000000000000000000000000111111010111111010111111011111111100111111110000000000000000000000000000;
        // mem[106] = 128'b00000000000000000000000000000000000000000000000000000000111100011111111000111010110111100101111111011000000000000000000000000000;
        // mem[107] = 128'b00000000000000000000000000000000000000000000000000000000111010110111010100111011010111010111111010110000000000000000000000000000;
        // mem[108] = 128'b00000000000000000000000000000000000000000000000000000000111011101111011000111100100111011110111011010000000000000000000000000000;
        // mem[109] = 128'b00000000000000000000000000000000000000000000000000000000111101100111100011111110100111101101111100100000000000000000000000000000;
        // mem[110] = 128'b00000000000000000000000000000000000000000000000000000000111110110111110100111111100111110101111110100000000000000000000000000000;
        // mem[111] = 128'b00000000000000000000000000000000000000000000000000000000111111010111111011111111011111111100111111100000000000000000000000000000;
        // mem[112] = 128'b00000000000000000000000000000000000000000000000000000000111111100111111011111111000111111011111111011000000000000000000000000000;
        // mem[113] = 128'b00000000000000000000000000000000000000000000000000000000111110100111111011111100111111110010111111000000000000000000000000000000;
        // mem[114] = 128'b00000000000000000000000000000000000000000000000000000000111100011111101001111100110111100010111100111000000000000000000000000000;
        // mem[115] = 128'b00000000000000000000000000000000000000000000000000000000111100100111100010111101011111101010111100110000000000000000000000000000;
        // mem[116] = 128'b00000000000000000000000000000000000000000000000000000000111100000111100011111011111111100111111101011000000000000000000000000000;
        // mem[117] = 128'b00000000000000000000000000000000000000000000000000000000111011001111011101111010110111011000111011111000000000000000000000000000;
        // mem[118] = 128'b00000000000000000000000000000000000000000000000000000000111010110111010110111010110111010101111010110000000000000000000000000000;
        // mem[119] = 128'b00000000000000000000000000000000000000000000000000000000111010110111010110111011000111011000111010110000000000000000000000000000;
        // mem[120] = 128'b00000000000000000000000000000000000000000000000000000000000001101000000000000001110000001110000000000000010000000010000000000000;
        // mem[121] = 128'b00000000000000000000000000000000000000000000000000000000000010001000001110000010010000001110000001110000010001000001111000010000;
        // mem[122] = 128'b00000000000000000000000000000000000000000000000000000000000011010000010110000011001000010110000010010000010101000010010000010001;
        // mem[123] = 128'b00000000000000000000000000000000000000000000000000000000000011101000011100000011010000011001000011001000010101000010100000010101;
        // mem[124] = 128'b00000000000000000000000000000000000000000000000000000000000100000000011110000011100000011100000011010000010111000010110000010101;
        // mem[125] = 128'b00000000000000000000000000000000000000000000000000000000000100010000100001000011110000011110000011100000011010000011001000010111;
        // mem[126] = 128'b00000000000000000000000000000000000000000000000000000000000100000000100001000100000000011111000011110000011011000011010000011010;
        // mem[127] = 128'b00000000000000000000000000000000000000000000000000000000000011110000100010000011100000011111000100000000011010000011100000011011;
        // mem[128] = 128'b00000000000000000000000000000000000000000000000000000000000011010000011100000011000000011100000011100000011010000011100000011010;
        // mem[129] = 128'b00000000000000000000000000000000000000000000000000000000000011000000011000000011001000011000000011000000011010000011001000011010;
        // mem[130] = 128'b00000000000000000000000000000000000000000000000000000000000011001000011001000010110000010110000011001000011000000010110000011010;
        // mem[131] = 128'b00000000000000000000000000000000000000000000000000000000000010111000011000000010101000010110000010110000010101000010110000011000;
        // mem[132] = 128'b00000000000000000000000000000000000000000000000000000000000010111000010110000011000000010110000010101000011001000010110000010101;
        // mem[133] = 128'b00000000000000000000000000000000000000000000000000000000000010111000010111000011100000011000000011000000011100000011011000011001;
        // mem[134] = 128'b00000000000000000000000000000000000000000000000000000000000011000000011010000011001000011010000011100000011001000011011000011100;
        // mem[135] = 128'b00000000000000000000000000000000000000000000000000000000000010110000010110000011000000010111000011001000011000000011000000011001;
        // mem[136] = 128'b00000000000000000000000000000000000000000000000000000000000010110000010101000010110000010110000011000000010111000011001000011000;
        // mem[137] = 128'b00000000000000000000000000000000000000000000000000000000000010101000010100000010010000010110000010110000010000000010110000010111;
        // mem[138] = 128'b00000000000000000000000000000000000000000000000000000000000001010000010011111111110000001010000010010111111101000000111000010000;
        // mem[139] = 128'b00000000000000000000000000000000000000000000000000000000111111001111111111111110110111111000111111110111110111111110111111111101;
        // mem[140] = 128'b00000000000000000000000000000000000000000000000000000000111110010111110100111110001111110000111110110111110010111110001111110111;
        // mem[141] = 128'b00000000000000000000000000000000000000000000000000000000111110100111110001111111011111110101111110001111111100111110110111110010;
        // mem[142] = 128'b00000000000000000000000000000000000000000000000000000000111111010111111000111110101111111011111111011111110111111111011111111100;
        // mem[143] = 128'b00000000000000000000000000000000000000000000000000000000111111001111110110111111001111110110111110101111111000111110111111110111;
        // mem[144] = 128'b00000000000000000000000000000000000000000000000000000000111111001111111100111110111111110111111111001111110101111110111111111000;
        // mem[145] = 128'b00000000000000000000000000000000000000000000000000000000111111010111111001111111001111111000111110111111110111111111000111110101;
        // mem[146] = 128'b00000000000000000000000000000000000000000000000000000000111110101111111001111110000111110110111111001111101111111110100111110111;
        // mem[147] = 128'b00000000000000000000000000000000000000000000000000000000111101011111110000111101010111101011111110000111101000111101011111101111;
        // mem[148] = 128'b00000000000000000000000000000000000000000000000000000000111101100111101011111101011111101011111101010111101011111101001111101000;
        // mem[149] = 128'b00000000000000000000000000000000000000000000000000000000111101011111101010111101011111101100111101011111101011111101100111101011;
        // mem[150] = 128'b00000000000000000000000000000000000000000000000000000000111101000111101010111101010111101001111101011111101010111101010111101011;
        // mem[151] = 128'b00000000000000000000000000000000000000000000000000000000111100110111101000111100101111100111111101010111101000111101001111101010;
        // mem[152] = 128'b00000000000000000000000000000000000000000000000000000000111100110111100100111101000111100101111100101111100111111100011111101000;
        // mem[153] = 128'b00000000000000000000000000000000000000000000000000000000111101001111101000111101001111101000111101000111101001111101000111100111;
        // mem[154] = 128'b00000000000000000000000000000000000000000000000000000000111101011111101001111101100111101010111101001111101001111101001111101001;
        // mem[155] = 128'b00000000000000000000000000000000000000000000000000000000111101011111101011111100111111101001111101100111101000111101001111101001;
        // mem[156] = 128'b00000000000000000000000000000000000000000000000000000000111100111111100111111101000111101000111100111111101010111101000111101000;
        // mem[157] = 128'b00000000000000000000000000000000000000000000000000000000111100101111100110111100000111100101111101000111100011111100110111101010;
        // mem[158] = 128'b00000000000000000000000000000000000000000000000000000000111011111111100001111011101111011111111100000111011100111100010111100011;
        // mem[159] = 128'b00000000000000000000000000000000000000000000000000000000111011100111011110111011100111011100111011101111011100111011101111011100;
        // mem[160] = 128'b00000000000000000000000000000000000000000000000000000000111011111111011110111100010111011111111011100111100010111011110111011100;
        // mem[161] = 128'b00000000000000000000000000000000000000000000000000000000111100101111100001111100111111100111111100010111101001111100111111100010;
        // mem[162] = 128'b00000000000000000000000000000000000000000000000000000000111101000111100111111101000111100110111100111111101000111101010111101001;
        // mem[163] = 128'b00000000000000000000000000000000000000000000000000000000111101000111100111111101100111101001111101000111101111111101001111101000;
        // mem[164] = 128'b00000000000000000000000000000000000000000000000000000000111101011111101101111100101111101010111101100111100101111101100111101111;
        // mem[165] = 128'b00000000000000000000000000000000000000000000000000000000111011110111100111111011011111011011111100101111011011111011101111100101;
        // mem[166] = 128'b00000000000000000000000000000000000000000000000000000000111011110111011100111011110111011110111011011111011110111011110111011011;
        // mem[167] = 128'b00000000000000000000000000000000000000000000000000000000111011011111011110111010111111011010111011110111010110111011010111011110;
        // mem[168] = 128'b00000000000000000000000000000000000000000000000000000000111010100111010110111010111111010101111010111111010110111010101111010110;
        // mem[169] = 128'b00000000000000000000000000000000000000000000000000000000111011000111010101111011000111011000111010111111010111111010111111010110;
        // mem[170] = 128'b00000000000000000000000000000000000000000000000000000000111011001111010111111011100111011001111011000111011100111011001111010111;
        // mem[171] = 128'b00000000000000000000000000000000000000000000000000000000111100001111011110111100111111100000111011100111100110111100001111011100;
        // mem[172] = 128'b00000000000000000000000000000000000000000000000000000000111100111111101001111101000111100110111100111111100101111100101111100110;
        // mem[173] = 128'b00000000000000000000000000000000000000000000000000000000111100100111101011111100111111100101111101000111100111111100101111100101;
        // mem[174] = 128'b00000000000000000000000000000000000000000000000000000000111101010111100101111110011111101011111100111111110011111101011111100111;
        // mem[175] = 128'b00000000000000000000000000000000000000000000000000000000111110011111110010111110000111110010111110011111110000111110010111110011;
        // mem[176] = 128'b00000000000000000000000000000000000000000000000000000000111101101111110001111101010111101101111110000111101010111101100111110000;
        // mem[177] = 128'b00000000000000000000000000000000000000000000000000000000111101100111101011111110000111101011111101010111110000111101100111101010;
        // mem[178] = 128'b00000000000000000000000000000000000000000000000000000000111110100111110010111110001111110010111110000111110010111110000111110000;
        // mem[179] = 128'b00000000000000000000000000000000000000000000000000000000111101110111110010111101100111101101111110001111101100111101110111110010;
        // mem[180] = 128'b00000000000000000000000000000000000000000000000000000000111101110111101011111110011111101111111101100111110010111101111111101100;
        // mem[181] = 128'b00000000000000000000000000000000000000000000000000000000111110010111110010111110010111110110111110011111110011111110011111110010;
        // mem[182] = 128'b00000000000000000000000000000000000000000000000000000000111101110111110000111101101111101110111110010111101100111101111111110011;
        // mem[183] = 128'b00000000000000000000000000000000000000000000000000000000111101011111101100111101101111101100111101101111101100111101011111101100;
        // mem[184] = 128'b00000000000000000000000000000000000000000000000000000000111110000111101100111110100111110001111101101111110101111110001111101100;
        // mem[185] = 128'b00000000000000000000000000000000000000000000000000000000111110101111110100111110011111110110111110100111110011111111000111110101;
        // mem[186] = 128'b00000000000000000000000000000000000000000000000000000000111101111111110011111101011111101110111110011111101011111101101111110011;
        // mem[187] = 128'b00000000000000000000000000000000000000000000000000000000111101101111101100111110010111101100111101011111110010111101101111101011;
        // mem[188] = 128'b00000000000000000000000000000000000000000000000000000000111111000111110010111111001111111000111110010111110111111111000111110010;
        // mem[189] = 128'b00000000000000000000000000000000000000000000000000000000111110100111111001111101111111110100111111001111110000111110100111110111;
        // mem[190] = 128'b00000000000000000000000000000000000000000000000000000000111110000111110000111110010111110000111101111111110010111101110111110000;
        // mem[191] = 128'b00000000000000000000000000000000000000000000000000000000111110010111110011111101110111110011111110010111101101111110010111110010;
        // mem[192] = 128'b00000000000000000000000000000000000000000000000000000000111101111111101111111111111111110010111101110111111110111101111111101101;
        // mem[193] = 128'b00000000000000000000000000000000000000000000000000000000000001010111111011000010000000001010111111111000001110000001011111111110;
        // mem[194] = 128'b00000000000000000000000000000000000000000000000000000000000011001000010101000010001000010100000010000000001100000001010000001110;
        // mem[195] = 128'b00000000000000000000000000000000000000000000000000000000000010010000010101000010010000010001000010001000001111000001110000001100;
        // mem[196] = 128'b00000000000000000000000000000000000000000000000000000000000010101000010100000010110000010100000010010000010011000010010000001111;
        // mem[197] = 128'b00000000000000000000000000000000000000000000000000000000000010111000010110000010110000010101000010110000010011000010011000010011;
        // mem[198] = 128'b00000000000000000000000000000000000000000000000000000000000010110000010110000010100000010101000010110000010101000010101000010011;
        // mem[199] = 128'b00000000000000000000000000000000000000000000000000000000000010101000010101000010100000010101000010100000010010000010011000010101;
        // mem[200] = 128'b00000000000000000000000000000000000000000000000000000000000010001000010001000010001000010011000010100000010001000010001000010010;
        // mem[201] = 128'b00000000000000000000000000000000000000000000000000000000000010010000010001000001111000001100000010001000001011000001101000010001;
        // mem[202] = 128'b00000000000000000000000000000000000000000000000000000000000011001000010110000011100000010110000001111000010011000010000000001011;
        // mem[203] = 128'b00000000000000000000000000000000000000000000000000000000000110110000100111000101011000100110000011100000011011000010110000010011;
        // mem[204] = 128'b00000000000000000000000000000000000000000000000000000000000111010000111010000110101000101111000101011000100010000011100000011011;
        // mem[205] = 128'b00000000000000000000000000000000000000000000000000000000000110110000111011000110110000111001000110101000111010000101111000100010;
        // mem[206] = 128'b00000000000000000000000000000000000000000000000000000000000010111000100100000100001000101100000110110000110001000111001000111010;
        // mem[207] = 128'b00000000000000000000000000000000000000000000000000000000000010101000010100000010100000010110000100001000011111000100111000110001;
        // mem[208] = 128'b00000000000000000000000000000000000000000000000000000000000010111000010101000010101000010110000010100000010101000011010000011111;
        // mem[209] = 128'b00000000000000000000000000000000000000000000000000000000000010101000010110000010011000010011000010101000010001000010011000010101;
        // mem[210] = 128'b00000000000000000000000000000000000000000000000000000000000010110000010101000010101000010101000010011000010001000010001000010001;
        // mem[211] = 128'b00000000000000000000000000000000000000000000000000000000000010001000010100000010000000010011000010101000001110000010001000010001;
        // mem[212] = 128'b00000000000000000000000000000000000000000000000000000000000010010000010000000010001000010000000010000000001101000001101000001110;
        // mem[213] = 128'b00000000000000000000000000000000000000000000000000000000000010100000010101000010011000010010000010001000001111000001100000001101;
        // mem[214] = 128'b00000000000000000000000000000000000000000000000000000000000010001000010011000010001000010100000010011000010100000010011000001111;
        // mem[215] = 128'b00000000000000000000000000000000000000000000000000000000000001001000001101000000001000001011000010001000000101000010000000010100;
        // mem[216] = 128'b00000000000000000000000000000000000000000000000000000000111111111000000010111111000111111101000000001111111010111111101000000101;
        // mem[217] = 128'b00000000000000000000000000000000000000000000000000000000111101100111111001111110000111110110111111000111111000111111010111111010;
        // mem[218] = 128'b00000000000000000000000000000000000000000000000000000000111011100111100111111010100111011111111110000111010100111100011111111000;
        // mem[219] = 128'b00000000000000000000000000000000000000000000000000000000111010111111010101111011000111010101111010100111011000111010110111010100;
        // mem[220] = 128'b00000000000000000000000000000000000000000000000000000000111011111111011000111100100111011110111011000111100011111011101111011000;
        // mem[221] = 128'b00000000000000000000000000000000000000000000000000000000111100111111100010111110000111101001111100100111110100111101100111100011;
        // mem[222] = 128'b00000000000000000000000000000000000000000000000000000000111110100111101110111111010111110100111110000111111011111110110111110100;
        // mem[223] = 128'b00000000000000000000000000000000000000000000000000000000111111100111110110111111101111111011111111010111111011111111010111111011;
        // mem[224] = 128'b00000000000000000000000000000000000000000000000000000000111111000111111011111111011111111011111111101111111011111111100111111011;
        // mem[225] = 128'b00000000000000000000000000000000000000000000000000000000111110001111110101111101100111110100111111011111101001111110100111111011;
        // mem[226] = 128'b00000000000000000000000000000000000000000000000000000000111100000111101000111100000111100011111101100111100010111100011111101001;
        // mem[227] = 128'b00000000000000000000000000000000000000000000000000000000111011101111011101111011110111011110111100000111100011111100100111100010;
        // mem[228] = 128'b00000000000000000000000000000000000000000000000000000000111101000111100001111011110111100010111011110111011101111100000111100011;
        // mem[229] = 128'b00000000000000000000000000000000000000000000000000000000111011101111100111111011000111011101111011110111010110111011001111011101;
        // mem[230] = 128'b00000000000000000000000000000000000000000000000000000000111011011111011001111011000111011000111011000111010110111010110111010110;
        // mem[231] = 128'b00000000000000000000000000000000000000000000000000000000111011001111011010111011000111011000111011000111011000111010110111010110;
        // mem[232] = 128'b00000000000000000000000000000000000000000000000000000000000010101000000000000010010000010001000000000000001110000001101000000000;
        // mem[233] = 128'b00000000000000000000000000000000000000000000000000000000000011011000010110000011010000010110000010010000010110000010001000001110;
        // mem[234] = 128'b00000000000000000000000000000000000000000000000000000000000011111000011110000011101000011100000011010000011100000011010000010110;
        // mem[235] = 128'b00000000000000000000000000000000000000000000000000000000000011111000011110000100000000011111000011101000011110000011101000011100;
        // mem[236] = 128'b00000000000000000000000000000000000000000000000000000000000100001000100000000100010000100001000100000000100001000100000000011110;
        // mem[237] = 128'b00000000000000000000000000000000000000000000000000000000000100001000100001000100100000100010000100010000100001000100010000100001;
        // mem[238] = 128'b00000000000000000000000000000000000000000000000000000000000100001000100010000100001000100001000100100000100010000100000000100001;
        // mem[239] = 128'b00000000000000000000000000000000000000000000000000000000000011110000100000000011101000100000000100001000011100000011110000100010;
        // mem[240] = 128'b00000000000000000000000000000000000000000000000000000000000011011000011011000011001000011010000011101000011000000011010000011100;
        // mem[241] = 128'b00000000000000000000000000000000000000000000000000000000000011000000011010000011000000011000000011001000011001000011000000011000;
        // mem[242] = 128'b00000000000000000000000000000000000000000000000000000000000011000000010110000011001000011001000011000000011000000011001000011001;
        // mem[243] = 128'b00000000000000000000000000000000000000000000000000000000000011010000010111000010111000011000000011001000010110000010111000011000;
        // mem[244] = 128'b00000000000000000000000000000000000000000000000000000000000011011000011011000011000000011001000010111000010111000010111000010110;
        // mem[245] = 128'b00000000000000000000000000000000000000000000000000000000000011010000011000000011001000011001000011000000011010000010111000010111;
        // mem[246] = 128'b00000000000000000000000000000000000000000000000000000000000010110000011000000010101000010111000011001000010110000011000000011010;
        // mem[247] = 128'b00000000000000000000000000000000000000000000000000000000000010011000010100000010011000010101000010101000010101000010110000010110;
        // mem[248] = 128'b00000000000000000000000000000000000000000000000000000000000010100000010100000010110000010100000010011000010100000010110000010101;
        // mem[249] = 128'b00000000000000000000000000000000000000000000000000000000000010011000010110000010001000010011000010110000010011000010101000010100;
        // mem[250] = 128'b00000000000000000000000000000000000000000000000000000000000001001000010001111111110000001000000010001111111111000001010000010011;
        // mem[251] = 128'b00000000000000000000000000000000000000000000000000000000111110111111111101111110011111111001111111110111110100111111001111111111;
        // mem[252] = 128'b00000000000000000000000000000000000000000000000000000000111110001111110110111110001111110001111110011111110001111110010111110100;
        // mem[253] = 128'b00000000000000000000000000000000000000000000000000000000111110111111110010111111011111110111111110001111111000111110100111110001;
        // mem[254] = 128'b00000000000000000000000000000000000000000000000000000000111111101111111101111111001111111100111111011111110110111111010111111000;
        // mem[255] = 128'b00000000000000000000000000000000000000000000000000000000111111100111111100111111111111111100111111001111111100111111001111110110;
        // mem[256] = 128'b00000000000000000000000000000000000000000000000000000000111111101000000000111111001111111100111111111111111001111111001111111100;
        // mem[257] = 128'b00000000000000000000000000000000000000000000000000000000111110110111111000111110111111111000111111001111111001111111010111111001;
        // mem[258] = 128'b00000000000000000000000000000000000000000000000000000000111110011111110110111101110111110100111110111111110000111110101111111001;
        // mem[259] = 128'b00000000000000000000000000000000000000000000000000000000111101010111101101111101010111101001111101110111101011111101011111110000;
        // mem[260] = 128'b00000000000000000000000000000000000000000000000000000000111101010111101010111101010111101011111101010111101010111101100111101011;
    end

    // read_pointer pointer
    always@(posedge m00_axis_aclk)
    begin
        if(!m00_axis_aresetn)
        begin
            read_pointer <= 0;
        end
        else if(send_tx)
        begin
            read_pointer <= read_pointer + 1'b1;
        end
        else
        begin
            read_pointer <= read_pointer;
        end
    end

    // stall counter increase
    always@(posedge m00_axis_aclk)
    begin
        if(!m00_axis_aresetn)
        begin
            stall_cnt <= 0;
        end
        else if(read_pointer >= (OUTPUT_WORD_ID_STALL_FOR_50_CYCLE - 1))
        begin
            stall_cnt <= stall_cnt + 1'b1;
        end
        else
        begin
            stall_cnt <= stall_cnt;
        end
    end

    always@(posedge m00_axis_aclk)
    begin
        if(!m00_axis_aresetn)
        begin
            m00_axis_tvalid_inner <= 1'b1;
        end
        else if (read_pointer == (OUTPUT_WORD_ID_STALL_FOR_50_CYCLE-1) && (stall_cnt < 50))
        begin
            m00_axis_tvalid_inner <= 1'b0;
        end
        else if (read_pointer == (OUTPUT_WORD_ID_STALL_FOR_50_CYCLE) && (stall_cnt >= 50))
        begin    
            m00_axis_tvalid_inner <= 1'b1;
        end
        else if(read_pointer == (NUMBER_OF_OUTPUT_WORDS-1))
        begin
            m00_axis_tvalid_inner <= 1'b0;
        end
        else
        begin
            m00_axis_tvalid_inner <= m00_axis_tvalid_inner;
        end
    end

    // read_pointer pointer
    always@(posedge m00_axis_aclk)
    begin
        if(!m00_axis_aresetn)
        begin
            no_send <= 1'b0;
        end
        else if (read_pointer == (OUTPUT_WORD_ID_STALL_FOR_50_CYCLE - 1) && (stall_cnt < 50))
        begin    
            no_send <= 1'b1;
        end
        else if (read_pointer == (OUTPUT_WORD_ID_STALL_FOR_50_CYCLE) && (stall_cnt >= 50))
        begin    
            no_send <= 1'b0;
        end
        else if (read_pointer == (NUMBER_OF_OUTPUT_WORDS-1))
        begin    
            no_send <= 1'b1;
        end
        else
        begin
            no_send <= no_send;
        end
    end

    // always@(posedge m00_axis_aclk)
    // begin
    //     if(!m00_axis_aresetn)
    //     begin
    //         m00_axis_tvalid_inner <= 1'b1;
    //     end
    //     else if(read_pointer == (NUMBER_OF_OUTPUT_WORDS-1))
    //     begin
    //         m00_axis_tvalid_inner <= 1'b0;
    //     end
    //     else
    //     begin
    //         m00_axis_tvalid_inner <= m00_axis_tvalid_inner;
    //     end
    // end

    // //read_pointer pointer
    // always@(posedge m00_axis_aclk)
    // begin
    //     if(!m00_axis_aresetn)
    //     begin
    //         no_send <= 1'b0;
    //     end
    //     else if (read_pointer == (NUMBER_OF_OUTPUT_WORDS-1))
    //     begin    
    //         no_send <= 1'b1;
    //     end
    //     else
    //     begin
    //         no_send <= no_send;
    //     end
    // end

    // read_pointer pointer
    always@(*)
    begin
        if(!m00_axis_aresetn)
        begin
            tx_done <= 1'b0;
        end
        else if (read_pointer == (NUMBER_OF_OUTPUT_WORDS-1))
        begin    
            tx_done <= 1'b1;
        end
        else
        begin
            tx_done <= 1'b0;
        end
    end

    // Streaming output data is read from FIFO
    always @(*)
    begin
        if(!m00_axis_aresetn)
        begin
            m00_axis_tdata_inner <= mem[0];
        end
        else if(no_send)
        begin
            m00_axis_tdata_inner <= 0;
        end
        else
        begin
            m00_axis_tdata_inner <= mem[read_pointer]; //read_pointer + 32'b1;
        end
    end

    assign  m00_axis_tvalid = m00_axis_tvalid_inner;
    assign  m00_axis_tdata = m00_axis_tdata_inner;
    assign  m00_axis_tstrb = {(C_M_AXIS_TDATA_WIDTH/8){m00_axis_tvalid_inner}};
    assign  m00_axis_tlast = tx_done;

endmodule
